module main

#flag -I @VMODROOT/src/c/
#flag @VMODROOT/src/c/tmp.o
#include "tmp.h"

fn C.test_func(voidptr, &char)
